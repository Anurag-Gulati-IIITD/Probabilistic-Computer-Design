module tanh_LUT(
    input [6 : 0] bias,
    output reg [31 : 0] tanh_out
);


    always @(*) begin
        case(bias) 
            7'b1100000: tanh_out = 32'b1_0000000000000000000000111100101;
            7'b1011111: tanh_out = 32'b1_0000000000000000000001100011110;
            7'b1011110: tanh_out = 32'b1_0000000000000000000010100100011;
            7'b1011101: tanh_out = 32'b1_0000000000000000000100001111000;
            7'b1011100: tanh_out = 32'b1_0000000000000000000110111110101;
            7'b1011011: tanh_out = 32'b1_0000000000000000001011100000010;
            7'b1011010: tanh_out = 32'b1_0000000000000000010010111101110;
            7'b1011001: tanh_out = 32'b1_0000000000000000011111010000111;
            7'b1011000: tanh_out = 32'b1_0000000000000000110011100010111;
            7'b1010111: tanh_out = 32'b1_0000000000000001010100111110101;
            7'b1010110: tanh_out = 32'b1_0000000000000010001100000110110;
            7'b1010101: tanh_out = 32'b1_0000000000000011100110111111010;
            7'b1010100: tanh_out = 32'b1_0000000000000101111100110101000;
            7'b1010011: tanh_out = 32'b1_0000000000001001110011110111000;
            7'b1010010: tanh_out = 32'b1_0000000000010000001011000111001;
            7'b1010001: tanh_out = 32'b1_0000000000011010101010011110010;
            7'b1010000: tanh_out = 32'b1_0000000000101011111101000111111;
            7'b1001111: tanh_out = 32'b1_0000000001001000011101000011000;
            7'b1001110: tanh_out = 32'b1_0000000001110111011010011101001;
            7'b1001101: tanh_out = 32'b1_0000000011000100110000110101010;
            7'b1001100: tanh_out = 32'b1_0000000101000100000101110111101;
            7'b1001011: tanh_out = 32'b1_0000001000010101011110110010110;
            7'b1001010: tanh_out = 32'b1_0000001101101101001111101101001;
            7'b1001001: tanh_out = 32'b1_0000010110100000000101001010001;
            7'b1001000: tanh_out = 32'b1_0000100100110101011111010001001;
            7'b1000111: tanh_out = 32'b1_0000111100000010000000110100010;
            7'b1000110: tanh_out = 32'b1_0001100001001000001101000100000;
            7'b1000101: tanh_out = 32'b1_0010011011010110111000100010100;
            7'b1000100: tanh_out = 32'b1_0011110100001000001010100101101;
            7'b1000011: tanh_out = 32'b1_0101110101100110111000001101100;
            7'b1000010: tanh_out = 32'b1_1000100110110010101100001010010;
            7'b1000001: tanh_out = 32'b1_1100000101001101000000101011010;
            7'b0000000: tanh_out = 32'b0_0000000000000000000000000000000;
            7'b0000001: tanh_out = 32'b0_0011111010110010111111010100110;
            7'b0000010: tanh_out = 32'b0_0111011001001101010011110101110;
            7'b0000011: tanh_out = 32'b0_1010001010011001000111110010100;
            7'b0000100: tanh_out = 32'b0_1100001011110111110101011010011;
            7'b0000101: tanh_out = 32'b0_1101100100101001000111011101100;
            7'b0000110: tanh_out = 32'b0_1110011110110111110010111100000;
            7'b0000111: tanh_out = 32'b0_1111000011111101111111001011110;
            7'b0001000: tanh_out = 32'b0_1111011011001010100000101110111;
            7'b0001001: tanh_out = 32'b0_1111101001011111111010110101111;
            7'b0001010: tanh_out = 32'b0_1111110010010010110000010010111;
            7'b0001011: tanh_out = 32'b0_1111110111101010100001001101010;
            7'b0001100: tanh_out = 32'b0_1111111010111011111010001000011;
            7'b0001101: tanh_out = 32'b0_1111111100111011001111001010110;
            7'b0001110: tanh_out = 32'b0_1111111110001000100101100010111;
            7'b0001111: tanh_out = 32'b0_1111111110110111100010111101000;
            7'b0010000: tanh_out = 32'b0_1111111111010100000010111000001;
            7'b0010001: tanh_out = 32'b0_1111111111100101010101100001110;
            7'b0010010: tanh_out = 32'b0_1111111111101111110100111000111;
            7'b0010011: tanh_out = 32'b0_1111111111110110001100001001000;
            7'b0010100: tanh_out = 32'b0_1111111111111010000011001011000;
            7'b0010101: tanh_out = 32'b0_1111111111111100011001000000110;
            7'b0010110: tanh_out = 32'b0_1111111111111101110011111001010;
            7'b0010111: tanh_out = 32'b0_1111111111111110101011000001011;
            7'b0011000: tanh_out = 32'b0_1111111111111111001100011101001;
            7'b0011001: tanh_out = 32'b0_1111111111111111100000101111001;
            7'b0011010: tanh_out = 32'b0_1111111111111111101101000010010;
            7'b0011011: tanh_out = 32'b0_1111111111111111110100011111110;
            7'b0011100: tanh_out = 32'b0_1111111111111111111001000001011;
            7'b0011101: tanh_out = 32'b0_1111111111111111111011110001000;
            7'b0011110: tanh_out = 32'b0_1111111111111111111101011011101;
            7'b0011111: tanh_out = 32'b0_1111111111111111111110011100010;
            7'b0100000: tanh_out = 32'b0_1111111111111111111111000011011;

            default: tanh_out = 32'b0;
        endcase
    end

endmodule