module tanh_LUT(
    input [5 : 0] bias,
    output reg [31 : 0] tanh_out
);


    always @(*) begin
        case(bias) 
            6'b111100: tanh_out = 32'b1_0000000000101011111101000111111;
            6'b111101: tanh_out = 32'b1_0000000101000100000101110111101;
            6'b111110: tanh_out = 32'b1_0000100100110101011111010001001;
            6'b111111: tanh_out = 32'b1_0011110100001000001010100101101;
            6'b000000: tanh_out = 32'b0_0000000000000000000000000000000;
            6'b000001: tanh_out = 32'b0_1100001011110111110101011010011;
            6'b000010: tanh_out = 32'b0_1111011011001010100000101110111;
            6'b000011: tanh_out = 32'b0_1111111010111011111010001000011;
            6'b000100: tanh_out = 32'b0_1111111111010100000010111000001;
            default: tanh_out = 32'b0;
        endcase
    end
    // always @(*) begin
    //     case(bias)
    //         6'b110000: tanh_out = 32'b1_111_1111_1110_1010_0000_0101_1100_0001;
    //         6'b110001: tanh_out = 32'b1_1111111110110111100010111101000;
    //         6'b110010: tanh_out = 32'b1_1111111110001000100101100010111;
    //         6'b110011: tanh_out = 32'b1_1111111100111011001111001010110;
    //         6'b110100: tanh_out = 32'b1_1111111010111011111010001000011;
    //         6'b110101: tanh_out = 32'b1_1111110111101010100001001101010;
    //         6'b110110: tanh_out = 32'b1_1111110010010010110000010010111;
    //         6'b110111: tanh_out = 32'b1_1111101001011111111010110101111;
    //         6'b111000: tanh_out = 32'b1_1111011011001010100000101110111;
    //         6'b111001: tanh_out = 32'b1_1111000011111101111111001011110;
    //         6'b111010: tanh_out = 32'b1_1110011110110111110010111100000;
    //         6'b111011: tanh_out = 32'b1_1101100100101001000111011101100;
    //         6'b111100: tanh_out = 32'b1_1100001011110111110101011010011;
    //         6'b111101: tanh_out = 32'b1_1010001010011001000111110010100;
    //         6'b111110: tanh_out = 32'b1_0111011001001101010011110101110;
    //         6'b111111: tanh_out = 32'b1_0011111010110010111111010100110;
    //         6'b000000: tanh_out = 32'b0_0000000000000000000000000000000;
    //         6'b000001: tanh_out = 32'b0_0011111010110010111111010100110;
    //         6'b000010: tanh_out = 32'b0_0111011001001101010011110101110;
    //         6'b000011: tanh_out = 32'b0_1010001010011001000111110010100;
    //         6'b000100: tanh_out = 32'b0_1100001011110111110101011010011;
    //         6'b000101: tanh_out = 32'b0_1101100100101001000111011101100;
    //         6'b000110: tanh_out = 32'b0_1110011110110111110010111100000;
    //         6'b000111: tanh_out = 32'b0_1111000011111101111111001011110;
    //         6'b001000: tanh_out = 32'b0_1111011011001010100000101110111;
    //         6'b001001: tanh_out = 32'b0_1111101001011111111010110101111;
    //         6'b001010: tanh_out = 32'b0_1111110010010010110000010010111;
    //         6'b001011: tanh_out = 32'b0_1111110111101010100001001101010;
    //         6'b001100: tanh_out = 32'b0_1111111010111011111010001000011;
    //         6'b001101: tanh_out = 32'b0_1111111100111011001111001010110;
    //         6'b001110: tanh_out = 32'b0_1111111110001000100101100010111;
    //         6'b001111: tanh_out = 32'b0_1111111110110111100010111101000;
    //         default: tanh_out = 32'b0;
    //     endcase
    // end

endmodule